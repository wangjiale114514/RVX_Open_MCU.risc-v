`include "../Units/RVX_Info.v"

module Stage_ID (
    input wire clk,
    input wire rst,
    input wire flush,                    // 清空流水线信号
);
    
endmodule